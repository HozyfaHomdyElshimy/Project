


module DW02_multp( a, b, tc, out0, out1 );


// parameters
parameter a_width = 8;
parameter b_width = 8;
parameter out_width = 18;

`define npp ((a_width/2) + 2)         //6
`define xdim (a_width+b_width+1)      //17
`define bsxt (a_width+1)               //9

//-----------------------------------------------------------------------------
 //I/O decalarations
input [a_width-1 : 0]	a;
input [b_width-1 : 0]	b;
input			tc;
output [out_width-1:0]	out0, out1;



//-----------------------------------------------------------------------------
// synopsys translate_off

reg   [`xdim-1 : 0]       pp_array [0 : `npp-1];    //17...6
reg   [`xdim-1 : 0]      	 tmp_OUT0, tmp_OUT1;    //17
wire  [a_width+2 : 0]	               a_padded;     //11
wire  [`xdim-1 : 0]                    b_padded;     //17
wire  [`xdim-b_width-1 : 0]      	temp_padded;     //9
wire  			       a_sign, b_sign, out_sign;

//-----------------------------------------------------------------------------

  
  initial begin : parameter_check
    integer param_err_flg;

    param_err_flg = 0;
    
    
    if (a_width < 1) begin
      param_err_flg = 1;
      $display(
	"ERROR: %m :\n  Invalid value (%d) for parameter a_width (lower bound: 1)",
	a_width );
    end
    
    if (b_width < 1) begin
      param_err_flg = 1;
      $display(
	"ERROR: %m :\n  Invalid value (%d) for parameter b_width (lower bound: 1)",
	b_width );
    end
    
    if (out_width < (a_width+b_width+2)) begin
      param_err_flg = 1;
      $display(
	"ERROR: %m :\n  Invalid value (%d) for parameter out_width (lower bound: (a_width+b_width+2))",
	out_width );
    end
  
    if ( param_err_flg == 1) begin
      $display(
        "%m :\n  Simulation aborted due to invalid parameter value(s)");
      $finish;
    end

  end // parameter_check

//-----------------------------------------------------------------------------

  assign a_sign = tc & a[a_width-1];
  assign b_sign = tc & b[b_width-1];
  assign a_padded = {a_sign, a_sign, a, 1'b0};
  assign temp_padded = {`bsxt{b_sign}};
  assign b_padded = {temp_padded, b};

  always @ (a_padded or b_padded)
  begin : mk_pp_array
    reg [`xdim-1 : 0] temp_pp_array [0 : `npp-1];
    reg [`xdim-1 : 0] next_pp_array [0 : `npp-1];
    reg [`xdim+3 : 0] temp_pp;
    reg [`xdim-1 : 0] new_pp;
    reg [`xdim-1 : 0] tmp_pp_carry;
    reg [a_width+2 : 0] temp_a_padded;
    reg [2 : 0] temp_bitgroup;
    integer bit_pair, pp_count, i;

    temp_pp_array[0] = {`xdim{1'b0}};

    for (bit_pair=0 ; bit_pair < `npp-1 ; bit_pair = bit_pair+1)
    begin
      temp_a_padded = (a_padded >> (bit_pair*2));
      temp_bitgroup = temp_a_padded[2 : 0];

      case (temp_bitgroup)
        3'b000, 3'b111 :
          temp_pp = {`xdim{1'b0}};
        3'b001, 3'b010 :
          temp_pp = b_padded;
        3'b011 :
          temp_pp = b_padded << 1;
        3'b100 :
          temp_pp = (~(b_padded << 1) + 1);
        3'b101, 3'b110 :
          temp_pp =  ~b_padded + 1;
        default : temp_pp = {`xdim{1'b0}};
      endcase

      temp_pp = temp_pp << (2 * bit_pair);
      new_pp = temp_pp[`xdim-1 : 0];
      temp_pp_array[bit_pair+1] = new_pp;
    end
    pp_count = `npp;

    while (pp_count > 2)
    begin
      for (i=0 ; i < (pp_count/3) ; i = i+1)
      begin
        next_pp_array[i*2] = temp_pp_array[i*3] ^ temp_pp_array[i*3+1] ^ temp_pp_array[i*3+2];

        tmp_pp_carry = (temp_pp_array[i*3] & temp_pp_array[i*3+1]) |
                       (temp_pp_array[i*3+1] & temp_pp_array[i*3+2]) |
                       (temp_pp_array[i*3] & temp_pp_array[i*3+2]);

        next_pp_array[i*2+1] = tmp_pp_carry << 1;
      end

      if ((pp_count % 3) > 0)
      begin
        for (i=0 ; i < (pp_count % 3) ; i = i + 1)
        next_pp_array[2 * (pp_count/3) + i] = temp_pp_array[3 * (pp_count/3) + i];
      end

      for (i=0 ; i < `npp ; i = i + 1) 
        temp_pp_array[i] = next_pp_array[i];

      pp_count = pp_count - (pp_count/3);
    end

    tmp_OUT0 <= temp_pp_array[0];

    if (pp_count > 1)
      tmp_OUT1 <= temp_pp_array[1];
    else
      tmp_OUT1 <= {`xdim{1'b0}};
  end // mk_pp_array


  assign out_sign = tmp_OUT0[`xdim-1 ] | tmp_OUT1[`xdim-1];
  assign out0 = ((^(a ^ a) !== 1'b0) | (^(b ^ b) !== 1'b0) | (^(tc ^ tc) !== 1'b0)) ? {out_width{1'bx}} 
                : {{out_width-`xdim{1'b0}}, tmp_OUT0};
  assign out1 = ((^(a ^ a) !== 1'b0) | (^(b ^ b) !== 1'b0) | (^(tc ^ tc) !== 1'b0)) ? {out_width{1'bx}} 
                : {{out_width-`xdim{out_sign}}, tmp_OUT1};

// synopsys translate_on
endmodule



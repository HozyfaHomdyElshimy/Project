`timescale 1ns / 1ps
module FloatAdditionTB ();

reg [31:0] A,B;
wire [31:0] result;
wire Flag_ADD;
real  value;

  reg                    RST,  clk  ;
  reg                       EN ;

FloatingAddition F_Add (.CLK(clk),.RST(RST),.Flag_ADD(Flag_ADD),.EN(EN),.A(A),.B(B),.OUT_ADD(result));


initial  
begin
 $display("\t\t  Time a b result ");
 $monitor("%d %b %b %b ", $time , A, B, result); 
 
 //initial values
clk = 1'b0;
EN = 1'b1 ;

A = 32'b1_11111111_00000000000000000000000;  // -inf
B = 32'b0_10000000_10011001100110011001100;  // 3.2
#20

A = 32'b01000001101100100110011001100110; // 22.3
B = 32'b10111111000000000000000000000000;  // -0.5
#20

A = 32'b01000001011111001100110011001101; // 15.8
B = 32'b00111111101001100110011001100110;  // 1.3
#20

A = 32'b01000010011000000000000000000000; // 56
B = 32'b00000000000000000000000000000000;  // 0
#20
A = 32'b0_01111110_01010001111010111000010;  // 0.66
B = 32'b0_01111110_00000101000111101011100;  // 0.51
#20
A = 32'b1_10000001_10011001100110011001100;  // -6.4 
B = 32'b1_01111110_00000000000000000000000;  // -0.5
#20
A = 32'b0_10000001_10011001100110011001100;  // 6.4
B = 32'b1_01111110_00000000000000000000000;  // -0.5
#20
A = 32'b1_01111110_00000000000000000000000;  // -0.5
B = 32'b0_10000001_10011001100110011001100;  // 6.4
#20
A = 32'b10111111100000000000000000000000;  // -1
B = 32'b01000000000000000000000000000000;  // 2
end
always #20 clk = ~clk;
endmodule
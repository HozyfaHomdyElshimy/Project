`timescale 1ns / 1ps
module F_Division_TB ();
reg [31:0] A,B;
reg clk,RST;
reg                       EN ;
reg overflow, underflow, exception;
wire [31:0] result;
//real  value;
F_Division F_Div (
.A(A),
.B(B),
.RST(RST),
.clk(clk),
.EN(EN),
.overflow(overflow),
.underflow(underflow),
.exception(exception),
.result(result));

initial  
begin
 $display("\t\t  Time a b result ");
 $monitor("%d %b %b %b ", $time , A, B, result); 
 
 
 //initial values
clk = 1'b0;
EN = 1'b1 ;

A = 32'b01000001000111000000000000000000;  // 9.75
B = 32'b01000000100000000000000000000000;  // 4
#20


A = 32'b00000000000000000000000000000000;   // 0
B = 32'b01000001000111000000000000000000;  // 9.75
//#20 
//A = 32'b00111111101001100110011001100110;    // 1.3
//B = 32'b00000000000000000000000000000000;   // 0
#20
A = 32'b01111111100000000000000000000000;   // inf
B = 32'b01000001000111000000000000000000;  // 9.75
//#20 
//A = 32'b00111111101001100110011001100110;    // 1.3
//B = 32'b01111111100000000000000000000000;  // inf
#20

A = 32'b01000001101100100110011001100110; // 22.3
B = 32'b10111111000000000000000000000000;  // -0.5
#20

A = 32'b0_01111110_01010001111010111000010;  // 0.66
B = 32'b0_01111110_00000101000111101011100;  // 0.51
#20
A = 32'b1_10000001_10011001100110011001100;  // -6.4 
B = 32'b1_01111110_00000000000000000000000;  // -0.5
#20
A = 32'b0_10000001_10011001100110011001100;  // 6.4
B = 32'b1_01111110_00000000000000000000000;  // -0.5

end
always #5 clk = ~clk;
endmodule
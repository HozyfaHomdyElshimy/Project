`timescale 1ns / 1ps

module FloatingMultiplication 
(input [31:0]                     A,
input [31:0]                      B,                
input  wire                       CLK ,
input  wire                       RST ,
input  wire                       EN ,
output                 infinity, zero,                      
output reg  [31:0]            OUT_MUL ,
output reg                  Flag_Mul);
                                 
                               
                                 
reg [23:0] A_Mantissa;
reg [23:0] B_Mantissa;
reg [22:0] Mantissa;
reg [47:0] Temp_Mantissa;
reg [7:0] A_Exponent,B_Exponent,Temp_Exponent,diff_Exponent,Exponent;
reg A_sign,B_sign,Sign;
reg [32:0] Temp;
reg [6:0] exp_adjust;
wire expones, expzeros, sigzeros;

  assign expones = (&A[30:23])|(&B[30:23]);
  assign expzeros = (~|A[30:23])|(~|B[30:23]);
  assign sigzeros = (~|A[22:0])|(~|B[22:0]);

   
  assign infinity       =  expones      &  sigzeros ;
  assign zero           =  expzeros     &  sigzeros ;
  
  always @ (posedge CLK or negedge RST)
 begin 
   if (!RST)
     begin
      OUT_MUL <= 'b0 ;
      Flag_Mul <= 'b0 ;	
	 end
   else
     begin   
      
//always@(*)
//begin
if (EN)
    begin

  if(infinity)
    begin
     OUT_MUL =32'b0_11111111_00000000000000000000000; //return default nan
    end
      else if (zero)
    begin
      OUT_MUL =32'b0_00000000_00000000000000000000000;
    end
  else
    begin
A_Mantissa = {1'b1,A[22:0]};
A_Exponent = A[30:23];
A_sign = A[31];
  
B_Mantissa = {1'b1,B[22:0]};
B_Exponent = B[30:23];
B_sign = B[31];

Temp_Exponent = A_Exponent+B_Exponent-127;
Temp_Mantissa = A_Mantissa*B_Mantissa;
Mantissa = Temp_Mantissa[47] ? Temp_Mantissa[46:24] : Temp_Mantissa[45:23];
Exponent = Temp_Mantissa[47] ? Temp_Exponent+1'b1 : Temp_Exponent;
Sign = A_sign^B_sign;
OUT_MUL = {Sign,Exponent,Mantissa};
end
end
end
end

endmodule



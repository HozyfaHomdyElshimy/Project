`timescale 1ns / 1ps

module F_Division
                        (input [31:0]                      A,
                         input [31:0]                      B,
                         input                             clk,
                         input                             RST,
                         input  wire                       EN ,
                         output                       overflow,
                         output                       underflow,
                         output                       exception,
                         output reg [31:0]              result);
                         
reg [23:0] A_Mantissa,B_Mantissa;
reg [22:0] Mantissa;
wire [7:0] exp;
reg [23:0] Temp_Mantissa;
reg [7:0] A_Exponent,B_Exponent,Temp_Exponent,diff_Exponent;
wire [7:0] Exponent;
reg [7:0] A_adjust,B_adjust;
reg A_sign,B_sign,Sign;
reg [32:0] Temp;
wire [31:0] temp1,temp2,temp3,temp4,temp5,temp6,temp7,debug;
wire [31:0] reciprocal;
wire [31:0] x0,x1,x2,x3;
reg [6:0] exp_adjust;
reg [31:0] B_scaled; 
reg en1,en2,en3,en4,en5;
reg dummy;
wire [31:0] result1;
wire    infinity, zero, MUL_enable,ADD_enable;


/*----Initial value----*/
F_Mul M1        //verified
(
.A({1'b0,8'd126,B[22:0]}),
.B(32'h3ff0f0f1),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_MUL(temp1),
.infinity(infinity),
.zero(zero)
);

assign debug = {1'b1,temp1[30:0]};
F_Addition A1
(
.A(32'h4034b4b5),
.B({1'b1,temp1[30:0]}),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_ADD(x0)
); 

/*----First Iteration----*/
F_Mul M2
(
.A({1'b0,8'd126,B[22:0]}),
.B(x0),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_MUL(temp2),
.infinity(infinity),
.zero(zero)
);

F_Addition A2
(
.A(32'h40000000),
.B({!temp2[31],temp2[30:0]}),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_ADD(temp3)
); 

F_Mul M3
(
.A(x0),
.B(temp3),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_MUL(x1),
.infinity(infinity),
.zero(zero)
);

/*----Second Iteration----*/
F_Mul M4
(
.A({1'b0,8'd126,B[22:0]}),
.B(x1),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_MUL(temp4),
.infinity(infinity),
.zero(zero)
);


F_Addition A3
(
.A(32'h40000000),
.B({!temp4[31],temp4[30:0]}),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_ADD(temp5)
); 

F_Mul M5
(
.A(x1),
.B(temp5),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_MUL(x2),
.infinity(infinity),
.zero(zero)
);


/*----Third Iteration----*/
F_Mul M6
(
.A({1'b0,8'd126,B[22:0]}),
.B(x2),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_MUL(temp6),
.infinity(infinity),
.zero(zero)
);

F_Addition A4
(
.A(32'h4034b4b5),
.B({1'b1,temp1[30:0]}),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_ADD(temp7)
); 

F_Mul M7
(
.A(x2),
.B(temp7),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_MUL(x3),
.infinity(infinity),
.zero(zero)
);

/*----Reciprocal : 1/B----*/
assign Exponent = x3[30:23]+8'd126-B[30:23];
assign reciprocal = {B[31],Exponent,x3[22:0]};

/*----Multiplication A*1/B----*/
F_Mul M8
(
.A(A),
.B(reciprocal),
.RST(RST),
.CLK(clk),
.EN(EN),
.OUT_MUL(result1),
.infinity(infinity),
.zero(zero)
);


always @(posedge clk or negedge RST)
begin
if (!EN || !RST)
    begin
      
      result  <= 'b0 ;
      	
	 end
   else
     begin
       result = result1;
     end
     end

endmodule